interface interf;
  logic clk;
  logic rst;
  logic en;
  logic [3:0]count;
endinterface
