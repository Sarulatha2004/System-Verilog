

rrgerg
