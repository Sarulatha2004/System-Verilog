module task_example;
  
  task compare(input int a,b, output done);
    if(a>b)
      $display("a is greater than b");
    else if(a <b)
      $display("a is less than b");
    else
      $display("a is equal to b");
    
    #10;
    done =1;
  endtask
  
  initial begin
    bit done;
    
    compare(10,10,done);
    if(done)
      $display("Comparison completed at a time=%0t",$time);
    compare(5,9,done);
    if(done)
      $display("Comparison completed at a time=%0t",$time);
    compare(9,5,done);
    if(done)
      $display("Comparison completed at a time=%0t",$time);
  end
endmodule
