interface fifo_inf #(parameter DATA_WIDTH=8);
  
  logic wclk;
  logic rclk;
  logic wrstn;
  logic rrstn;
  logic r_en;
  logic w_en;
  logic [DATA_WIDTH-1:0]data_in;
  logic [DATA_WIDTH-1:0]data_out;
  logic full;
  logic empty;
  
endinterface
  
  
