module fifo_mem #(parameter DEPTH=8, DATA_WIDTH=8,PTR_WIDTH=3)
  
  (
    input logic wclk,
    input logic rclk,
    input logic w_en,
    input logic r_en,
    input logic [PTR_WIDTH:0]b_wptr,
    input logic [PTR_WIDTH:0]b_rptr,
    input logic [DATA_WIDTH-1:0]data_in,
    input logic full,
    input logic empty,
    output logic [DATA_WIDTH-1:0]data_out
  );
  
  
  logic [DATA_WIDTH-1:0]fifo [DEPTH-1:0];
  
  
  always_ff @(posedge wclk) begin
    
    if(w_en & !full)
      fifo[b_wptr[PTR_WIDTH-1:0]] <=data_in;
  end
  
  always_ff @(posedge rclk) begin
    
    if(r_en & !empty)
      data_out <= fifo[b_rptr[PTR_WIDTH-1:0]];
  end
  
  
endmodule
      
  
