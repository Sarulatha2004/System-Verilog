 module cons_repeat_bin;

  bit [3:0] a;
   bit [2:0] values[$] = '{2,6,2,8,2,2,4,4,4};

  covergroup cvgrp;
    c1 : coverpoint a {
      bins tran_1 = (2 [*2]);
      bins tran_2 = (4 [*3]); 
    }
  endgroup

  cvgrp cg = new();

  initial
  begin
    foreach(values[i])
    begin
      a = values[i];
      cg.sample();
      $display("val = %d, cov = %.2f %%", a, cg.get_inst_coverage());
    end
  end
endmodule


////////////OUTPUT/////////////////////


# KERNEL: val =  2, cov = 0.00 %
# KERNEL: val =  6, cov = 0.00 %
# KERNEL: val =  2, cov = 0.00 %
# KERNEL: val =  0, cov = 0.00 %
# KERNEL: val =  2, cov = 0.00 %
# KERNEL: val =  2, cov = 50.00 %
# KERNEL: val =  4, cov = 50.00 %
# KERNEL: val =  4, cov = 50.00 %
# KERNEL: val =  4, cov = 100.00 %

///////////////////////////////////////////
